interface xgemac_clk_interface();
  logic clk;
endinterface
