interface xgemac_rst_interface(input clk);
  logic rst;
endinterface
